//-----------------------------------------------------------------------------
//
// Title       : VDS_TB
// Design      : VehicleDetectSystem
// Author      : Kjersti
// Company     : NTNU
//
//-----------------------------------------------------------------------------
//
// File        : c:\My_Designs\VehicleDetectSystem\VehicleDetectSystem\src\VDS_TB.v
// Generated   : Mon Nov 21 12:39:21 2016
// From        : interface description file
// By          : Itf2Vhdl ver. 1.22
//
//-----------------------------------------------------------------------------
//
// Description : Testbench for complete digital part of Vehicle Detect System
//
//-----------------------------------------------------------------------------
`timescale 1 ns / 1 ns

//{{ Section below this comment is automatically maintained
//   and may be overwritten
//{module {VDS_TB}}
module VDS_TB ();  
	//Inputs to system
	reg fm0; //Data sent to decoder
	reg reset; //Reset signal for decoder and listener
	reg clk_50MHz; //50MHz clock for FSM in listener
	
	//System outputs
	wire interrupt;	//Interrupt signal from listener
	wire clk_500kHz; //Clock generated by decoder
	wire nrz; //NRZ signal from decoder
	
	reg clk_fm0; //Clock for timing input of FM0 signal
	
	//Message components:
	parameter flag		= 8'b01111110;
	parameter address 	= 8'b11111111; 
	parameter mac 		= 8'b10000000;
	parameter llc		= 8'b00000011;
	parameter infoT		= 8'b01010101; //Info when Emergency Vehicle nearby
	parameter infoF		= 8'b00110110; //Random info (no emergency vehicle)
	parameter FCST		= 16'b0010111111111010; //Correct FCS field when infoT
	parameter FCSF		= 16'b0011011110010010;	//Random (wrong) FCS field
	parameter preamble  = 8'b01010101;	
	
	//Message components added together to make complete message sequences:
	parameter infoN 	= {flag, address, mac, llc, infoF, FCST, flag}; //No emergency vehicle, wrong FCS
	parameter infoEV 	= {flag, address, mac, llc, infoT, FCST, flag};	//Emergency vehicle, right FCS
	parameter wrongFCS 	= {flag, address, mac, llc, infoT, FCSF, flag};	//Emergency vehicle, wrong FCS
	
	integer count;  
	reg [447:0] fm0_msg; //Holds FM0 test sequence
	reg [2:0] outputTB; //Signal used during simulation to show which information is being sent
	
	//Possible values of outputTB signal
	parameter s0_reset = 3'b000, s1_preamble = 3'b001, s2_infoN = 3'b010, s3_infoEV = 3'b011, s4_wrongFCS = 3'b100;
	
	//Declaration of test modules
	decoder decoderTest (.fm0(fm0), .reset(reset), .clk(clk_500kHz), .nrz(nrz));
	listener listenerTest (.nrz(nrz), .reset(reset), .clk_50MHz(clk_50MHz), .clk_500kHz(clk_500kHz), .interrupt(interrupt));
	
	//Function to convert 224 bit data(nrz) sequence to 448 bit FM0 sequence:
	function [447:0] bitsToFM0;
		input [223:0] nrzBits; //224 bit nrz sequence
		integer i;
		begin
			for(i = 447; i >= 0; i = i - 2) begin
				if(i == 447)
					bitsToFM0[i] = 1'b1;
				else
					bitsToFM0[i] = !bitsToFM0[i+1];
				
				if(nrzBits[(i-1)/2] == 1'b1)
					bitsToFM0[i-1] = bitsToFM0[i];
				else
					bitsToFM0[i-1] = !bitsToFM0[i];	
			end
		end
	endfunction
	
		
	//Initial setup
	initial 
		begin
			clk_50MHz = 0;
			clk_fm0 = 0;
			reset = 1;
			//Create FM0 input-sequence
			fm0_msg = bitsToFM0({preamble, infoN, preamble, infoEV, preamble, wrongFCS, preamble});
			////Content of fm0_msg: [447:432]preamble, [431:304]infoN, [303:288]preamble, [287:160]infoEV,  
			////[159:144]preamble, [143:16]wrongFCS, [15:0]preamble
			#1000
			reset = 0;
		end
		
	always @(posedge clk_fm0) begin
		if(reset == 1) //Reset
			begin
			fm0 = 1'b0;
			count = 447; //To be used as index when sending FM0 sequence 
			outputTB <= s0_reset;
			end
		else 
			begin
			fm0 = fm0_msg[count]; //Output FM0 sequence serially
			count = count - 1; //Index of fm0_msg
			//Change outputTB to show which part of fm0_msg is being sent:
			if((count > 303) && (count < 432))
				outputTB <= s2_infoN;
			else if((count > 159) && (count < 288))
				outputTB <= s3_infoEV;
			else if((count > 15) && (count < 144))
				outputTB <= s4_wrongFCS;
			else
				outputTB <= s1_preamble;
			end
	end 
	
	
	always begin//Clock generation, 50MHz clock
		#10 clk_50MHz = !clk_50MHz;
	end	
	
	always begin //Clock generation, FM0 clock for sending FM0 signal
		#500 clk_fm0 = !clk_fm0;
	end
	
endmodule
